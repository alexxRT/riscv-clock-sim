module testbench();

    reg clk = 1'b0;
    wire[31:0] WriteData;
    wire[31:0] DataAdr;
    reg reset;

    // instantiate device to be tested
    top testdevice(.clk(clk),      .WriteDataM(WriteData),
                   .reset(reset),  .ALUResultM(DataAdr)
    );

    // initialize test
    initial begin
        reset = 1; #17; reset = 0;
    end

    // generate clock to sequence tests
    always begin
        clk <= ~clk; #5;
    end


    initial begin
        $dumpvars;
        $display("Test started...");
        #1000
        $finish;
    end


endmodule